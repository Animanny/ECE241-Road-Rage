module drawBackground(input clk, reset, enable, output[7:0] x, output [6:0] y, output [2:0] colour);
		backgroundImage bG(.address(memCounter),.clock(clk),.q(colour));//iterate through address and read colour from memory
		
	//assign ledr = memCounter;
	
	reg[14:0] memCounter;// = 10'b1;
	reg[7:0] xCounter;// = 8'b0;
	reg[6:0] yCounter;// = 8'b0;
	initial begin
		memCounter = 10'b0;
		xCounter = 8'b0;
		yCounter = 7'b0;
	end
		
	always@(posedge clk) begin
		if(reset == 1)begin
			xCounter <= 8'b0;
			yCounter <= 7'b0;
			memCounter <= 15'b0;
		end
		else if(enable)begin
			if (memCounter < 15'd19200) begin
				if(xCounter < 8'd159)begin
					xCounter <= xCounter +  1'b1;
				end
				else begin
					xCounter <= 0;
					yCounter <= yCounter + 1'b1;
				end
				memCounter <= memCounter + 1'b1;
			end
			else begin
				xCounter <= 8'b0;
				yCounter <= 7'b0;
				memCounter <= 15'b0;
			end
		end
	end
	
	assign x = xCounter;
	assign y = yCounter;

endmodule

