//module vga_demo(CLOCK_50, SW, KEY,
//				VGA_R, VGA_G, VGA_B,
//				VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_CLK);
//	
//	input CLOCK_50;
//	input [17:0] SW;
//	input [1:0] KEY;
//	output [9:0] VGA_R;
//	output [9:0] VGA_G;
//	output [9:0] VGA_B;
//	output VGA_HS;
//	output VGA_VS;
//	output VGA_BLANK;
//	output VGA_SYNC;
//	output VGA_CLK;				
//
//	vga_adapter VGA(
//			.resetn(KEY[0]),
//			.clock(CLOCK_50),
//			.colour(SW[17:15]),
//			.x(SW[14:7]),
//			.y(SW[6:0]),
//			.plot(~(KEY[1])),
//			/* Signals for the DAC to drive the monitor. */
//			.VGA_R(VGA_R),
//			.VGA_G(VGA_G),
//			.VGA_B(VGA_B),
//			.VGA_HS(VGA_HS),
//			.VGA_VS(VGA_VS),
//			.VGA_BLANK(VGA_BLANK),
//			.VGA_SYNC(VGA_SYNC),
//			.VGA_CLK(VGA_CLK));
//		defparam VGA.RESOLUTION = "160x120";
//		defparam VGA.MONOCHROME = "FALSE";
//		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
//		defparam VGA.BACKGROUND_IMAGE = "crappy road.mif";
//		
//endmodule